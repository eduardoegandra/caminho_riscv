// Módulo para instrução LB
module lb_operation(
    input [31:0] mem_data,
    output [31:0] result
);
    assign result = mem_data;
endmodule
